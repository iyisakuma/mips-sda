LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY datapath IS
  PORT (
    clock, reset : IN std_logic;

    -- sinais de controle
    RegDst, RegWrite, ALUSrc : IN std_logic;
    MemWrite, MemToReg      : IN std_logic;
    ALUCtrl                 : IN std_logic_vector(2 downto 0);
	 Jump                    : IN std_logic;
	 PC_jump                 : IN std_logic_vector(9 downto 0);
    -- instrução (para PC)
    instruction_out         : OUT std_logic_vector(31 downto 0)
  );
END datapath;

ARCHITECTURE arc OF datapath IS

  COMPONENT arithmetic_logic_unit
    PORT (
      sel : IN  std_logic_vector(2 downto 0);
      A,B : IN  std_logic_vector(31 downto 0);
      F   : OUT std_logic_vector(31 downto 0)
    );
  END COMPONENT;

  COMPONENT register_file
    PORT (
      load_enable, clock, reset : IN std_logic;
      data                      : IN std_logic_vector(31 downto 0);
      destination_select        : IN std_logic_vector(3 downto 0);
      A_select, B_select        : IN std_logic_vector(3 downto 0);
      A_data, B_data            : OUT std_logic_vector(31 downto 0)
    );
  END COMPONENT;

  COMPONENT instructions_memory
    PORT (
      clock        : IN  std_logic;
      write_enable : IN  std_logic;
      write_address: IN  std_logic_vector(9 downto 0);
      read_address : IN  std_logic_vector(9 downto 0);
      data_in      : IN  std_logic_vector(31 downto 0);
      data_out     : OUT std_logic_vector(31 downto 0)
    );
  END COMPONENT;

  COMPONENT data_memory
    PORT (
      clock        : IN  std_logic;
      write_enable : IN  std_logic;
      write_address: IN  std_logic_vector(9 downto 0);
      read_address : IN  std_logic_vector(9 downto 0);
      data_in      : IN  std_logic_vector(31 downto 0);
      data_out     : OUT std_logic_vector(31 downto 0)
    );
  END COMPONENT;

  COMPONENT mux2_1
    GENERIC (N : INTEGER := 32);
    PORT (
      sel     : IN  std_logic;
      X0, X1  : IN  std_logic_vector(N-1 downto 0);
      out_mux : OUT std_logic_vector(N-1 downto 0)
    );
  END COMPONENT;

  -- sinais internos
  SIGNAL PC, PC_JUMP             : std_logic_vector(9 downto 0) := (others=>'0');
  SIGNAL instr           : std_logic_vector(31 downto 0);
  SIGNAL regA, regB      : std_logic_vector(31 downto 0);
  SIGNAL aluB, aluOut    : std_logic_vector(31 downto 0);
  SIGNAL memOut, wbData  : std_logic_vector(31 downto 0);
  SIGNAL destReg         : std_logic_vector(4 downto 0);
  SIGNAL imm_ext         : std_logic_vector(31 downto 0);

BEGIN

  -- PC
  PROCESS(clock)
  BEGIN
  IF rising_edge(clock) THEN
     IF Jump = '1' THEN
      PC <= PC_jump;
     ELSE
		PC <= std_logic_vector(unsigned(PC) + 1);
     END IF;
	 END IF;
	END PROCESS;

  -- Instruction memory
  imem: instructions_memory
    PORT MAP (
      clock => clock,
      write_enable => '0',
      write_address => (others=>'0'),
      read_address => PC,
      data_in => (others=>'0'),
      data_out => instr
    );

  instruction_out <= instr;

  -- Sign extend imediato
  imm_ext <= (31 downto 16 => instr(15)) & instr(15 downto 0);

  -- RegDst MUX
  mux_rd: mux2_1
    GENERIC MAP (N=>5)
    PORT MAP (
      sel => RegDst,
      X0  => instr(20 downto 16),
      X1  => instr(15 downto 11),
      out_mux => destReg
    );

  -- Register File
  regs: register_file
    PORT MAP (
      load_enable => RegWrite,
      clock => clock,
      reset => reset,
      data => wbData,
      destination_select => destReg(3 downto 0),
      A_select => instr(25 downto 21),
      B_select => instr(20 downto 16),
      A_data => regA,
      B_data => regB
    );

  -- ALUSrc MUX
  mux_alu: mux2_1
    PORT MAP (
      sel => ALUSrc,
      X0  => regB,
      X1  => imm_ext,
      out_mux => aluB
    );

  -- ALU
  alu: arithmetic_logic_unit
    PORT MAP (
      sel => ALUCtrl,
      A => regA,
      B => aluB,
      F => aluOut
    );

  -- Data memory
  dmem: data_memory
    PORT MAP (
      clock => clock,
      write_enable => MemWrite,
      write_address => aluOut(9 downto 0),
      read_address  => aluOut(9 downto 0),
      data_in => regB,
      data_out => memOut
    );

  -- MemToReg MUX
  mux_wb: mux2_1
    PORT MAP (
      sel => MemToReg,
      X0  => aluOut,
      X1  => memOut,
      out_mux => wbData
    );

END arc;
