library verilog;
use verilog.vl_types.all;
entity mips_vlg_vec_tst is
end mips_vlg_vec_tst;
